** Profile: "SCHEMATIC1-Resposta freq�encial"  [ C:\Users\j.mendez.orero\Desktop\Practica1\practica1-pspicefiles\schematic1\resposta freq�encial.sim ] 

** Creating circuit file "Resposta freq�encial.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Cadence\SPB_16.5\tools\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 50 1kHz 10MegHz
.PROBE V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
